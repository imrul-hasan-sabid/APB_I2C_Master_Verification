/*
+-------------------+---------+----------+---------+----------+---------+--------+--+------------------------+
| Operation         | arbitr  | start    | restart | sla_sent | write   | ack    |  |       status_code      |
|                   | _lost   |          |         |          |         |        |  +----+----+----+----+----+
|                   |         |          |         |          |         |        |  | Y4 | Y3 | Y2 | Y1 | Y0 |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| ARBITRATION_LOST  | 1       | x        | x       | x        | x       | x      |  |  0 | 0  | 1  | 1  | 1  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| START COMP        | 0       | 1        | x       | x        | x       | x      |  |  0 | 0  | 0  | 0  | 1  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| REP_START COMP    | 0       | 0        | 1       | x        | x       | x      |  |  0 | 0  | 0  | 1  | 0  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| SLA+W -> ACK      | 0       | 0        | 0       | 1        | 0       | 0      |  |  0 | 0  | 0  | 1  | 1  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| SLA+W -> NACK     | 0       | 0        | 0       | 1        | 0       | 1      |  |  0 | 0  | 1  | 0  | 0  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| SLA+R -> ACK      | 0       | 0        | 0       | 1        | 1       | 0      |  |  0 | 1  | 0  | 0  | 0  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| SLA+R -> NACK     | 0       | 0        | 0       | 1        | 1       | 1      |  |  0 | 1  | 0  | 0  | 1  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| DATA_SENT -> ACK  | 0       | 0        | 0       | 0        | 0       | 0      |  |  0 | 0  | 1  | 0  | 1  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| DATA_SENT -> NACK | 0       | 0        | 0       | 0        | 0       | 1      |  |  0 | 0  | 1  | 1  | 0  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| DATA_RCV -> ACK   | 0       | 0        | 0       | 0        | 1       | 0      |  |  0 | 1  | 0  | 1  | 0  |
+-------------------+---------+----------+---------+----------+---------+--------+  +----+----+----+----+----+
| DATA_RCV -> NACK  | 0       | 0        | 0       | 0        | 1       | 1      |  |  0 | 1  | 0  | 1  | 1  |
+-------------------+---------+----------+---------+----------+---------+--------+--+----+----+----+----+----+
*/



module  status_code_generator #(
        `include "twi_parameters.sv"
)(
        input   logic   sla_sent, 
        input   logic   write, 
        input   logic   ack_bit, 
        input   logic   start_en, 
        input   logic   restart_en, 
        input   logic   arbitration_lost,

        output  logic   [TWS_WIDTH-1:0] status_code_generator_status_value
); 

	assign status_code_generator_status_value[0] 	= arbitration_lost | start_en | ( ~restart_en & ~write & ~ack_bit) | (~restart_en & write & ack_bit); 
	assign status_code_generator_status_value[1] 	= arbitration_lost | (~start_en & (  restart_en | (~sla_sent & ack_bit) | (~sla_sent&write) | (sla_sent & ~write & ~ack_bit)    )) ;
	assign status_code_generator_status_value[2]	= arbitration_lost | (~start_en  & ~restart_en & ~write & (~sla_sent | ack_bit)); 
	assign status_code_generator_status_value[3]	= ~arbitration_lost & ~start_en & ~restart_en & write; 
        assign status_code_generator_status_value[4]    = 0; 
        
endmodule 
